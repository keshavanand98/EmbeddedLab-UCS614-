module hello;
initial begin
$display("hello World");
end
endmodule
